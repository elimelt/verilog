/* Testbench for Homework 3 Problem 1 */
module fifo_tb ();

	// for you to implement

	initial begin
	
		// for you to implement
		
	end  // initial
	
endmodule  // fifo_tb
